module q(b,e);
input [3:0]b;
output [3:0]e;



endmodule
module eighttoone(i,s,f);
input [7:0]i;
input [2:0]s;
output f;
reg f;
always @(i,s)
begin
	case(s)
	0:f=i[0];
	1:f=i[1];
	2:f=i[2];
	3:f=i[3];
	4:f=i[4];
	5:f=i[5];
	6:f=i[6];
	7:f=i[7];
	endcase
end
endmodule
