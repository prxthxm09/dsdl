module q(g,b);
input [3:0]g;
output [3:0]b;
always @(g)
begin

end
endmodule
